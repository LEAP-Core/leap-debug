typedef Bit#(32) MEM_DATA_SM;
typedef Bit#(14) MEM_ADDRESS;
typedef Bit#(14) WORKING_SET;
typedef Bit#(32) CYCLE_COUNTER;
typedef 3        N_SCRATCH;

