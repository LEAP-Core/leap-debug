`include "awb/provides/coh_mem_test_common.bsh"
typedef Bit#(64) CYCLE_COUNTER;

typedef `COH_MEM_TEST_ENGINE_NUM N_TOTAL_ENGINES;
typedef Bit#(TAdd#(TLog#(TAdd#(N_TOTAL_ENGINES,1)),1)) ENGINE_PORT_NUM;
typedef Bit#(`COH_MEM_TEST_MEMORY_ADDR_BITS) MEM_ADDRESS;
typedef Bit#(64) TEST_DATA;

`ifndef COH_MEM_TEST_DUAL_FPGA_ENABLE_Z
    typedef TDiv#(N_TOTAL_ENGINES,2) N_LOCAL_ENGINES;
`else
    typedef N_TOTAL_ENGINES N_LOCAL_ENGINES;
`endif
typedef TSub#(N_TOTAL_ENGINES, N_LOCAL_ENGINES) N_REMOTE_ENGINES;

typedef enum
{
    COH_TEST_REQ_WRITE_RAND,
    COH_TEST_REQ_WRITE_SEQ,
    COH_TEST_REQ_READ_RAND,
    COH_TEST_REQ_READ_SEQ,
    COH_TEST_REQ_RANDOM,
    COH_TEST_REQ_FENCE,
    COH_TEST_REQ_RANDOM_FENCE
}
COH_MEM_ENGINE_TEST_REQ
    deriving (Bits, Eq);

